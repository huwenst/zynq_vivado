`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/12/05 09:37:57
// Design Name: 
// Module Name: Divider
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Divider(
	input iClk100M,
	input iRstN,
	input [31:0]iA,
	input [31:0]iB,
	  input iEn,
	output [31:0]oS,
	output [31:0]oC,
	output oValida
    );

	
endmodule
